
module audio_mem();

endmodule 