
module pcm();

endmodule 